E8
07
00
20
6D
05
00
08
73
05
00
08
75
05
00
08
77
05
00
08
79
05
00
08
7B
05
00
08
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
7D
05
00
08
7F
05
00
08
00
00
00
00
81
05
00
08
83
05
00
08
85
05
00
08
85
05
00
08
85
05
00
08
85
05
00
08
85
05
00
08
85
05
00
08
85
05
00
08
85
05
00
08
85
05
00
08
85
05
00
08
85
05
00
08
85
05
00
08
85
05
00
08
85
05
00
08
9F
04
00
08
85
05
00
08
85
05
00
08
85
05
00
08
00
00
00
00
85
05
00
08
85
05
00
08
85
05
00
08
85
05
00
08
B9
04
00
08
D5
04
00
08
85
05
00
08
85
05
00
08
85
05
00
08
85
05
00
08
85
05
00
08
85
05
00
08
85
05
00
08
00
F0
02
F8
00
F0
3A
F8
0A
A0
90
E8
00
0C
82
44
83
44
AA
F1
01
07
DA
45
01
D1
00
F0
2F
F8
AF
F2
09
0E
BA
E8
0F
00
13
F0
01
0F
18
BF
FB
1A
43
F0
01
03
18
47
B0
0B
00
00
D0
0B
00
00
10
3A
24
BF
78
C8
78
C1
FA
D8
52
07
24
BF
30
C8
30
C1
44
BF
04
68
0C
60
70
47
00
00
00
23
00
24
00
25
00
26
10
3A
28
BF
78
C1
FB
D8
52
07
28
BF
30
C1
48
BF
0B
60
70
47
1F
B5
1F
BD
10
B5
10
BD
00
F0
37
FA
11
46
FF
F7
F7
FF
00
F0
55
F9
00
F0
55
FA
03
B4
FF
F7
F2
FF
03
BC
00
F0
59
FA
00
00
10
B5
01
20
55
49
88
60
00
BF
54
48
00
68
00
F0
04
00
04
28
F9
D1
02
20
50
49
C8
60
08
63
50
48
48
60
00
BF
4D
48
00
68
00
F0
02
00
02
28
F9
D1
4A
48
C0
69
40
F0
08
00
48
49
C8
61
18
20
49
49
08
60
46
48
C0
69
20
F0
08
00
44
49
C8
61
08
46
C0
68
40
F4
82
70
C8
60
00
BF
40
48
00
68
00
F0
08
00
08
28
F9
D1
3D
48
00
6B
40
F4
82
70
3B
49
08
63
00
F0
07
F9
00
F0
E6
F8
00
F0
DC
F8
00
F0
8F
F8
4F
F6
FF
70
38
49
08
60
34
48
C0
69
37
49
40
EA
01
00
31
49
C8
61
35
48
88
62
4F
F0
E0
60
48
62
10
BD
33
48
34
49
88
60
00
20
08
60
4F
F6
FF
70
C8
60
00
20
48
60
40
1E
88
61
00
06
2F
49
88
60
00
20
08
60
4F
F6
FF
70
C8
60
4F
F4
7F
40
48
60
4F
F0
FF
30
88
61
29
48
2A
49
88
60
00
20
08
60
4F
F6
FF
70
C8
60
46
F6
FF
10
48
60
4F
F0
FF
30
88
61
24
48
25
49
88
60
00
20
08
60
4F
F6
FF
70
C8
60
48
60
4F
F0
FF
30
88
61
20
48
21
49
88
60
4F
F6
FF
70
1D
49
C8
60
40
1E
48
60
4F
F0
FF
30
1C
49
88
61
70
47
02
20
1B
49
48
62
20
20
88
62
60
20
C8
62
40
F2
01
30
08
63
70
47
00
20
16
49
C8
60
08
60
42
F2
0F
70
48
60
09
20
88
60
02
20
88
65
01
20
C8
60
70
47
00
00
00
00
02
40
04
0B
B1
00
00
80
01
40
BC
00
00
30
00
C0
41
24
00
00
04
04
55
55
55
C1
00
80
0A
40
00
00
0B
40
55
55
FF
FF
00
80
0B
40
55
55
00
54
00
80
0C
40
5A
55
55
55
00
80
0E
40
00
00
0D
40
00
00
07
40
00
BF
3A
48
80
6B
10
F4
80
4F
FA
D0
70
47
70
B5
03
46
0E
46
03
B9
70
BD
02
B9
FC
E7
1C
46
34
48
31
18
00
25
06
E0
34
F8
02
0B
21
F8
02
0B
FF
F7
E7
FF
6D
1C
95
42
F6
D3
00
BF
EC
E7
70
B5
03
46
0E
46
03
B9
70
BD
02
B9
FC
E7
1C
46
06
F1
40
51
00
25
06
E0
34
F8
02
0B
21
F8
02
0B
FF
F7
D0
FF
6D
1C
95
42
F6
D3
00
BF
EC
E7
22
49
00
20
03
E0
00
22
21
F8
02
2B
40
1C
B0
F5
7F
4F
F8
D3
70
47
1B
49
00
20
03
E0
00
22
21
F8
02
2B
40
1C
B0
F5
80
3F
F8
D3
70
47
15
48
80
6B
4F
F6
FB
71
08
40
12
49
88
63
70
47
11
48
80
6B
4F
F6
FE
71
08
40
0E
49
88
63
70
47
0D
48
80
6B
48
F2
10
01
08
43
0A
49
88
63
08
46
80
6B
4F
F6
FD
71
08
40
07
49
88
63
70
47
05
48
80
6B
4F
F6
F7
71
08
40
03
49
88
63
70
47
0F
20
01
49
88
63
70
47
00
00
02
40
00
00
02
30
00
02
00
30
4F
F0
00
60
52
49
08
60
FF
F7
AE
FE
FF
F7
FE
FE
FF
F7
49
FF
FF
F7
3C
FF
FF
F7
AB
FF
FF
F7
B4
FF
00
24
0E
E0
4B
4B
03
EB
C4
03
5A
88
49
4B
33
F8
34
30
59
00
47
4B
03
EB
C4
03
58
68
FF
F7
82
FF
64
1C
04
2C
EE
D3
00
24
0E
E0
43
4B
03
EB
C4
03
5A
88
41
4B
33
F8
34
30
59
00
3F
4B
03
EB
C4
03
58
68
FF
F7
58
FF
64
1C
04
2C
EE
D3
FF
F7
B6
FF
FF
F7
A5
FF
18
20
01
21
81
40
42
09
4F
F0
E0
23
03
EB
82
02
C2
F8
00
11
00
BF
00
20
33
49
08
60
33
49
08
60
33
49
08
60
33
49
08
60
04
E0
2F
48
00
68
40
1C
2D
49
08
60
F9
E7
00
20
2F
49
48
65
2B
48
00
68
2E
49
08
60
29
48
00
68
40
1C
28
49
08
60
70
47
10
20
4F
F0
40
51
88
67
25
48
00
68
27
49
08
60
23
48
00
68
40
1C
22
49
08
60
70
47
01
20
4F
F0
40
51
88
67
1F
48
00
68
C0
02
20
49
08
60
1D
48
00
68
40
1C
1B
49
08
60
70
47
10
B5
0A
46
00
BF
1B
4B
9B
69
03
F0
80
03
80
2B
F9
D1
00
21
18
E0
03
88
C3
F3
07
23
16
4C
23
60
00
BF
14
4B
9B
69
03
F0
80
03
80
2B
F9
D1
10
F8
04
4B
E3
B2
10
4C
23
60
00
BF
0E
4B
9B
69
03
F0
80
03
80
2B
F9
D1
49
1C
91
42
E4
D3
10
BD
70
47
00
00
08
ED
00
E0
C4
00
00
20
00
00
00
20
B0
00
00
20
B4
00
00
20
B8
00
00
20
BC
00
00
20
00
00
07
40
00
00
0B
40
00
00
0D
40
09
48
09
48
00
47
FE
E7
FE
E7
FE
E7
FE
E7
FE
E7
FE
E7
FE
E7
FE
E7
FE
E7
FE
E7
00
00
03
48
04
49
04
4A
05
4B
70
47
00
00
C1
00
00
08
E8
01
00
20
E8
07
00
20
E8
03
00
20
E8
03
00
20
70
47
70
47
70
47
75
46
00
F0
28
F8
AE
46
05
00
69
46
53
46
20
F0
07
00
85
46
18
B0
20
B5
FF
F7
DF
FF
BD
E8
20
40
4F
F0
00
06
4F
F0
00
07
4F
F0
00
08
4F
F0
00
0B
21
F0
07
01
AC
46
AC
E8
C0
09
AC
E8
C0
09
AC
E8
C0
09
AC
E8
C0
09
8D
46
70
47
04
46
AF
F3
00
80
20
46
FF
F7
A5
FD
00
48
70
47
84
01
00
20
01
49
18
20
AB
BE
FE
E7
26
00
02
00
70
47
F8
76
7F
00
FF
FF
F8
76
7E
00
FF
FF
F8
76
7D
00
FF
FF
F8
76
7C
00
FF
FF
F8
76
7B
00
FF
FF
F8
76
7A
00
FF
FF
F8
76
77
00
FF
FF
F8
76
76
00
FF
FF
F8
76
73
00
FF
FF
F8
76
72
00
FF
FF
F8
76
6F
00
FF
FF
F8
76
6E
00
FF
FF
F8
76
6B
00
00
00
F8
76
6A
00
00
00
F8
76
67
00
00
00
F8
76
66
00
30
01
F8
76
65
00
00
00
F8
76
64
00
00
01
F8
76
63
00
00
00
F8
76
62
00
00
00
00
FC
FF
EE
95
F4
00
80
00
10
45
F8
2F
81
00
71
12
00
E2
76
04
00
00
00
00
71
12
00
E2
76
06
00
00
00
00
71
12
00
E2
76
04
00
02
00
00
71
12
00
E2
76
06
00
AD
00
00
71
12
00
E2
76
04
00
03
00
00
71
12
00
E2
76
06
00
00
00
00
71
12
00
E2
76
04
00
04
00
00
71
12
00
E2
76
06
00
AD
00
00
71
12
00
E2
76
04
00
05
00
00
71
12
00
E2
76
06
00
00
00
00
71
12
00
E2
76
04
00
06
00
00
71
12
00
E2
76
06
00
1F
00
00
71
12
00
E2
76
04
00
07
00
00
71
12
00
E2
76
06
00
4A
20
00
71
12
00
E2
76
04
00
09
00
00
71
12
00
E2
76
06
00
00
FF
00
71
12
00
E2
76
04
00
08
00
00
71
12
00
E2
76
06
00
00
FF
00
71
12
00
E2
76
04
00
0A
00
00
71
12
00
E2
76
06
00
FF
FF
00
71
12
00
E2
76
04
00
0B
00
00
71
12
00
E2
76
06
00
FF
FF
00
71
12
00
E2
76
04
00
0C
00
00
71
12
00
E2
76
06
00
FF
FF
00
71
12
00
E2
76
04
00
0D
00
00
71
12
00
E2
76
06
00
FF
FF
00
71
12
00
E2
76
04
00
0E
00
00
71
12
00
E2
76
06
00
00
3F
00
71
12
00
E2
76
04
00
01
00
00
71
12
00
E2
76
06
00
00
00
00
71
12
00
E2
76
04
00
00
00
00
71
12
00
E2
76
06
00
0F
01
01
EE
00
FC
FE
EE
95
F4
00
80
08
E8
00
6F
41
0D
03
F6
00
F0
00
01
01
80
20
F0
20
00
00
6F
03
0C
01
71
12
00
08
48
E2
4E
06
00
04
10
03
00
10
F0
01
00
01
71
12
00
08
48
E2
4E
04
00
B8
F6
01
10
00
F0
02
00
12
88
20
F0
FF
FC
82
18
40
F0
00
01
82
80
01
71
12
00
E2
69
02
00
00
0C
01
10
00
F0
02
00
12
88
20
F0
FF
CF
82
18
40
F0
00
10
82
80
01
10
00
F0
02
00
12
88
20
F0
FF
3F
82
18
40
F0
00
40
82
80
01
10
00
F0
03
00
12
88
20
F0
0F
C0
04
11
10
F3
01
00
30
F3
FF
03
E4
F3
82
18
A0
F1
82
81
01
10
00
F0
03
00
12
88
20
F0
F8
FF
82
18
40
F0
01
00
82
80
00
6F
41
0C
F8
32
08
00
02
E8
82
F4
F8
80
74
00
02
EE
00
FC
FD
EE
BB
F7
1D
77
88
FF
95
F4
95
F4
95
F4
F8
76
00
00
00
00
F8
76
01
00
FF
FF
F8
76
5E
00
FF
FF
F8
76
3C
00
00
00
F8
76
3D
00
00
00
95
F4
95
F4
F8
76
3A
00
FF
FF
F8
76
39
00
5F
09
F8
71
39
00
38
00
F8
76
3A
00
00
00
74
F2
89
80
20
F0
20
00
74
F2
89
80
20
F0
28
00
74
F2
89
80
20
F0
30
00
F8
76
3B
00
00
00
F8
69
00
00
08
00
F8
76
01
00
FF
FF
BB
F6
F8
76
85
01
3F
00
95
F4
F8
10
85
01
44
F8
D1
81
BB
F7
F8
76
85
01
3F
00
00
76
40
20
01
76
20
00
74
F2
00
80
20
F0
00
20
F8
76
3C
00
01
80
BB
F6
73
F0
D1
81
95
F4
08
4A
09
4A
0A
4A
12
4A
06
4A
07
4A
1D
4A
F8
68
07
00
3F
7D
F8
69
07
00
00
40
F8
68
1D
00
FC
FF
95
F4
F8
10
85
01
45
F8
01
82
F8
6B
85
01
FF
FF
95
F4
12
72
85
01
95
F4
E2
70
00
40
85
01
E2
70
00
20
85
01
1D
8A
07
8A
06
8A
12
8A
0A
8A
09
8A
08
8A
EB
F4
07
4A
1D
4A
F8
68
07
00
3F
7D
F8
69
07
00
00
40
F8
68
1D
00
FC
FF
95
F4
1D
8A
07
8A
9B
F4
11
4A
16
4A
FF
EE
F8
10
83
01
E3
F4
11
72
60
01
F8
10
11
00
45
F8
3A
82
11
48
00
F0
61
01
16
88
95
F4
95
F4
EE
10
FF
FF
E3
F4
E9
6C
FF
FF
34
82
F8
10
82
01
45
F8
41
82
F8
10
82
01
E3
F4
F8
10
81
01
45
F8
48
82
F8
10
81
01
E3
F4
F8
10
84
01
E3
F4
74
F0
71
82
73
F0
4D
82
11
4A
11
88
F8
10
83
01
E3
F4
B8
F7
20
E8
F8
08
60
01
46
F8
61
82
F8
10
84
01
E3
F4
73
F2
6F
82
95
F4
01
E8
12
72
60
01
12
48
00
F0
01
00
F8
80
60
01
E2
70
61
01
11
00
F8
10
84
01
E3
F4
00
E8
11
8A
00
FC
95
F4
73
F0
72
82
18
77
80
00
F8
6B
18
00
7F
00
F8
68
18
00
FE
FF
B8
F7
BE
F7
B9
F6
A0
F4
B7
F6
B5
F6
B6
F6
20
F0
3C
80
00
F1
01
00
4D
F8
A0
82
B8
F6
95
F4
20
F0
3C
80
73
F0
9A
82
F8
7E
12
00
00
F0
01
00
F8
47
11
00
92
7E
F8
00
11
00
00
F0
01
00
F8
7E
11
00
00
F0
01
00
89
6C
8F
82
B8
F7
FC
EE
20
F0
FF
FF
00
F1
01
00
4D
F8
B8
82
B8
F6
95
F4
20
F0
FF
FF
73
F2
B2
82
02
4E
95
F4
E3
F5
02
56
00
7E
00
11
4C
FA
B0
82
03
6B
01
00
B8
F6
04
EE
74
F0
94
81
74
F0
22
82
00
FC
F8
80
83
01
00
FC
F8
80
84
01
00
FC
01
00
60
01
00
00
01
00
81
01
00
00
01
00
82
01
00
00
01
00
83
01
BE
82
01
00
84
01
BE
82
00
00
06
4A
07
4A
FF
EE
B8
F7
B9
F7
BA
F4
B9
F4
13
88
04
71
12
00
05
10
10
88
10
F0
03
00
13
49
04
09
4D
FA
20
80
1A
88
95
F4
72
F2
1A
80
98
E5
58
E5
BB
6D
98
E5
58
E5
BB
6D
73
F2
35
80
98
E5
58
E5
BB
6D
EA
6D
02
00
72
F2
34
80
13
48
12
49
20
F6
42
FA
30
80
92
10
8A
11
98
E5
14
E5
8B
81
83
80
BB
6D
EA
6D
02
00
13
48
12
49
C0
F0
70
FD
01
E8
01
EE
07
8A
06
8A
00
FC
73
F2
94
81
18
77
00
01
EB
F6
95
F4
95
F4
95
F4
EB
F6
95
F4
95
F4
95
F4
EB
F6
95
F4
95
F4
95
F4
EB
F6
95
F4
95
F4
95
F4
EB
F6
95
F4
95
F4
95
F4
EB
F6
95
F4
95
F4
95
F4
EB
F6
95
F4
95
F4
95
F4
EB
F6
95
F4
95
F4
95
F4
EB
F6
95
F4
95
F4
95
F4
EB
F6
95
F4
95
F4
95
F4
EB
F6
95
F4
95
F4
95
F4
EB
F6
95
F4
95
F4
95
F4
EB
F6
95
F4
95
F4
95
F4
EB
F6
95
F4
95
F4
95
F4
EB
F6
95
F4
95
F4
95
F4
EB
F6
95
F4
95
F4
95
F4
EB
F6
95
F4
95
F4
95
F4
EB
F6
95
F4
95
F4
95
F4
73
F2
E8
81
95
F4
95
F4
73
F2
13
82
95
F4
95
F4
EB
F6
95
F4
95
F4
95
F4
73
F2
E8
81
95
F4
95
F4
EB
F6
95
F4
95
F4
95
F4
EB
F6
95
F4
95
F4
95
F4
73
F2
E8
81
95
F4
95
F4
EB
F6
95
F4
95
F4
95
F4
EB
F6
95
F4
95
F4
95
F4
EB
F6
95
F4
95
F4
95
F4
73
F2
13
82
95
F4
95
F4
EB
F6
95
F4
95
F4
95
F4
EB
F4
95
F4
01
00
00
00
C4
0C
00
08
00
00
00
20
C4
00
00
00
FC
00
00
08
88
0D
00
08
C4
00
00
20
24
07
00
00
18
01
00
08
4C
80
79
02
1A
06
00
08
3C
80
10
00
0C
0B
00
08
00
80
3C
00
2C
0B
00
08
80
FF
7E
00
A4
0B
00
08
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
40
00
00
30
50
00
00
30
60
00
00
30
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
