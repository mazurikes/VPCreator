@0	0800056D
@1	08000579
@2	00000000
@3	00000000
@4	08000585
@5	08000585
@6	08000585
@7	08000585
@8	08000585
@9	08000585
@A	08000585
@B	08000585
@C	F83AF000
@D	45DA0701
@E	F013000F
@F	00000BB0
@10	0752D8FA
@11	00004770
@12	D8FBC178
@13	BD1FB51F
@14	F000FFF7
@15	F000BC03
@16	4854BF00
@17	60C84950
@18	0002F000
@19	61C84948
@1A	49440008
@1B	4840BF00
@1C	F4406B00
@1D	F000F8E6
@1E	48346008
@1F	62884835
@20	20006088
@21	61881E40
@22	60C870FF
@23	492A4829
@24	10FFF646
@25	20006088
@26	618830FF
@27	1E4060C8
@28	491B2002
@29	63083001
@2A	6048700F
@2B	00004770
@2C	300000BC
@2D	400A8000
@2E	54005555
@2F	400D0000
@30	D0FA4F80
@31	E7FCB902
@32	F8210B02
@33	E7ECBF00
@34	461CE7FC
@35	0B02F821
@36	4922E7EC
@37	4F7FF5B0
@38	2B02F821
@39	F64F6B80
@3A	F64F6B80
@3B	F2486B80
@3C	71FDF64F
@3D	71F7F64F
@3E	47706388
@3F	6000F04F
@40	FF49F7FF
@41	E00E2400
@42	00593034
@43	2C041C64
@44	4B41885A
@45	F7FF6858
@46	FFA5F7FF
@47	0282EB03
@48	60084933
@49	1C406800
@4A	6800482B
@4B	47706008
@4C	60084927
@4D	F04F2001
@4E	481D6008
@4F	BF00460A
@50	E0182100
@51	699B4B14
@52	4C10B2E3
@53	D1F92B80
@54	E000ED08
@55	200000B4
@56	400B0000
@57	E7FEE7FE
@58	0000E7FE
@59	080000C1
@5A	200003E8
@5B	000546AE
@5C	F7FFB520
@5D	F04F0700
@5E	09C0E8AC
@5F	4770468D
@60	47704800
@61	00020026
@62	76F8FFFF
@63	FFFF007B
@64	007676F8
@65	76F8FFFF
@66	0000006B
@67	006676F8
@68	76F80100
@69	F495EEFF
@6A	000476E2
@6B	00127100
@6C	00AD0006
@6D	76E20012
@6E	71000004
@6F	000476E2
@70	00127100
@71	001F0006
@72	76E20012
@73	71000009
@74	000476E2
@75	00127100
@76	FFFF0006
@77	76E20012
@78	7100000C
@79	000476E2
@7A	00127100
@7B	3F000006
@7C	76E20012
@7D	71000000
@7E	F495EEFE
@7F	80010100
@80	4EE24808
@81	48080012
@82	F0208812
@83	69E20012
@84	CFFFF020
@85	88120002
@86	F0001001
@87	F3300001
@88	0003F000
@89	6F008082
@8A	EE020074
@8B	F495F495
@8C	005E76F8
@8D	F4950000
@8E	71F8095F
@8F	F0208089
@90	F0208089
@91	76F80008
@92	10F8F495
@93	7600003F
@94	76F82000
@95	4A094A08
@96	7D3F0007
@97	10F8F495
@98	7212F495
@99	01852000
@9A	F4EB8A08
@9B	40000007
@9C	4A11F49B
@9D	10F80160
@9E	F4958816
@9F	10F88234
@A0	018110F8
@A1	F4E30184
@A2	018310F8
@A3	10F88261
@A4	01607212
@A5	00110161
@A6	F073F495
@A7	001868F8
@A8	F6B6F6B5
@A9	F495F6B8
@AA	0001F000
@AB	7EF80001
@AC	F020EEFC
@AD	F020F495
@AE	7E005602
@AF	F074EE04
@B0	80F8FC00
@B1	00000181
@B2	01840001
@B3	F4BAF7B9
@B4	0003F010
@B5	801AF272
@B6	8035F273
@B7	48138034
@B8	E514E598
@B9	F0C04912
@BA	8194F273
@BB	F495F6EB
@BC	F495F6EB
@BD	F495F6EB
@BE	F495F6EB
@BF	F495F6EB
@C0	F495F6EB
@C1	F495F6EB
@C2	F495F6EB
@C3	F495F6EB
@C4	8213F273
@C5	81E8F273
@C6	F495F6EB
@C7	F495F6EB
@C8	F495F6EB
@C9	F495F6EB
@CA	08000CC4
@CB	08000D88
@CC	0279804C
@CD	003C8000
@CE	00000000
@CF	00000000
@D0	00000000
@D1	00000000
@D2	00000000
@D3	00000000
@D4	00000000
@D5	00000000
@D6	30000040
@D7	00000000
@D8	00000000
