@0	08000573
@1	0800057B
@2	00000000
@3	08000581
@4	08000585
@5	08000585
@6	08000585
@7	0800049F
@8	00000000
@9	08000585
@A	08000585
@B	08000585
@C	E890A00A
@D	F000D101
@E	BF180F01
@F	00000BD0
@10	C830BF24
@11	24002300
@12	BF280752
@13	BD10B510
@14	F000F955
@15	0000FA59
@16	F0006800
@17	48506308
@18	D1F92802
@19	49492018
@1A	460861C8
@1B	F0006800
@1C	493B7082
@1D	F000F8DC
@1E	493769C0
@1F	60E0F04F
@20	F64F6008
@21	492F0600
@22	407FF44F
@23	20006088
@24	F04F6048
@25	F64F6008
@26	49214820
@27	F04F6048
@28	20206248
@29	20004770
@2A	60882009
@2B	40020000
@2C	2441C000
@2D	400B0000
@2E	400C8000
@2F	40070000
@30	B5704770
@31	4834461C
@32	F7FF0B02
@33	4603B570
@34	5140F106
@35	FFD0F7FF
@36	E0032000
@37	4770D3F8
@38	F5B01C40
@39	400871FB
@3A	400871FE
@3B	43080110
@3C	49074008
@3D	49034008
@3E	40020000
@3F	60084952
@40	FF3CF7FF
@41	EB034B4B
@42	EB034B47
@43	2400D3EE
@44	3034F833
@45	1C64FF58
@46	21012018
@47	1100F8C2
@48	60084933
@49	6008492D
@4A	6008492E
@4B	F04F2010
@4C	68004823
@4D	67885140
@4E	1C406800
@4F	699B4B1B
@50	F3C38803
@51	0380F003
@52	BF006023
@53	42911C49
@54	200000C4
@55	200000B8
@56	400D0000
@57	E7FEE7FE
@58	49044803
@59	200001E8
@5A	47704770
@5B	46534669
@5C	E8BDFFDF
@5D	F04F0800
@5E	09C0E8AC
@5F	F3AF4604
@60	20000184
@61	76F84770
@62	FFFF007D
@63	007A76F8
@64	76F8FFFF
@65	FFFF006F
@66	006A76F8
@67	76F80130
@68	00000063
@69	10008000
@6A	71000000
@6B	000476E2
@6C	00127100
@6D	00000006
@6E	76E20012
@6F	71000005
@70	000476E2
@71	00127100
@72	204A0006
@73	76E20012
@74	71000008
@75	000476E2
@76	00127100
@77	FFFF0006
@78	76E20012
@79	7100000D
@7A	000476E2
@7B	00127100
@7C	00000006
@7D	76E20012
@7E	E8088000
@7F	0020F020
@80	10040006
@81	00044EE2
@82	1882FCFF
@83	0C000002
@84	F0401882
@85	3FFFF020
@86	88120003
@87	F3E403FF
@88	F0208812
@89	32F80C41
@8A	EEFDFC00
@8B	000076F8
@8C	76F8FFFF
@8D	76F8F495
@8E	00380039
@8F	F2740020
@90	76F80030
@91	FFFF0001
@92	F8440185
@93	76012040
@94	8001003C
@95	4A124A0A
@96	000769F8
@97	F8450185
@98	F4950185
@99	8A078A1D
@9A	4A1D4A07
@9B	001D68F8
@9C	EEFF4A16
@9D	F8450011
@9E	10EEF495
@9F	F8450182
@A0	8248F845
@A1	8271F074
@A2	F7B8F4E3
@A3	F4E30184
@A4	F0004812
@A5	018410F8
@A6	77188272
@A7	F7B8FFFE
@A8	803CF020
@A9	803CF020
@AA	001147F8
@AB	F0000011
@AC	F100FFFF
@AD	F273FFFF
@AE	FA4C1100
@AF	F0748194
@B0	FC000184
@B1	01820001
@B2	000082BE
@B3	8813F4B9
@B4	09044913
@B5	E558E598
@B6	E558E598
@B7	F6204912
@B8	8083818B
@B9	E801FD70
@BA	01007718
@BB	F495F495
@BC	F495F495
@BD	F495F495
@BE	F495F495
@BF	F495F495
@C0	F495F495
@C1	F495F495
@C2	F495F495
@C3	F495F495
@C4	F495F495
@C5	F495F495
@C6	F495F495
@C7	F495F495
@C8	F495F495
@C9	F495F495
@CA	20000000
@CB	200000C4
@CC	0800061A
@CD	08000B2C
@CE	00000000
@CF	00000000
@D0	00000000
@D1	00000000
@D2	00000000
@D3	00000000
@D4	00000000
@D5	00000000
@D6	30000050
@D7	00000000
@D8	00000000
