@0	08000575
@1	00000000
@2	0800057D
@3	08000583
@4	08000585
@5	08000585
@6	08000585
@7	08000585
@8	08000585
@9	080004B9
@A	08000585
@B	08000585
@C	44820C00
@D	F2AFF82F
@E	F0431AFB
@F	BF243A10
@10	BF44C130
@11	26002500
@12	BF48C130
@13	FA37F000
@14	B403FA55
@15	2001B510
@16	28040004
@17	BF006048
@18	69C0484A
@19	48466008
@1A	F44068C0
@1B	28080008
@1C	F0006308
@1D	F64FF88F
@1E	0001EA40
@1F	BD106248
@20	60C870FF
@21	20006088
@22	F04F6048
@23	F64F6008
@24	618830FF
@25	60C870FF
@26	F64F6088
@27	491C30FF
@28	20606288
@29	60C84916
@2A	65882002
@2B	00B10B04
@2C	04040000
@2D	FFFF5555
@2E	5555555A
@2F	483ABF00
@30	460E4603
@31	25001831
@32	1C6DFFE7
@33	B903460E
@34	E0062500
@35	42951C6D
@36	F8212200
@37	2000491B
@38	D3F83F80
@39	63884912
@3A	6388490E
@3B	6388490A
@3C	47706388
@3D	47706388
@3E	30020000
@3F	FEAEF7FF
@40	FFABF7FF
@41	885A03C4
@42	685803C4
@43	4B43E00E
@44	4B3F0059
@45	D3EE2C04
@46	09424081
@47	2000BF00
@48	60084933
@49	2000E7F9
@4A	68004829
@4B	67885140
@4C	49221C40
@4D	6800481F
@4E	6008491B
@4F	0380F003
@50	4C162307
@51	D1F92B80
@52	699B4B0E
@53	BD10D3E4
@54	20000000
@55	200000BC
@56	48094809
@57	E7FEE7FE
@58	4B054A04
@59	200007E8
@5A	46754770
@5B	0007F020
@5C	F04F4020
@5D	F0210B00
@5E	09C0E8AC
@5F	46208000
@60	20184901
@61	FFFF007F
@62	007C76F8
@63	76F8FFFF
@64	FFFF0073
@65	006E76F8
@66	76F80000
@67	00000065
@68	006276F8
@69	812FF845
@6A	76E20012
@6B	71000002
@6C	000476E2
@6D	00127100
@6E	00AD0006
@6F	76E20012
@70	71000006
@71	000476E2
@72	00127100
@73	FF000006
@74	76E20012
@75	7100000A
@76	000476E2
@77	00127100
@78	FFFF0006
@79	76E20012
@7A	7100000E
@7B	000476E2
@7C	00127100
@7D	010F0006
@7E	0D416F00
@7F	0C036F00
@80	F0100003
@81	1001F6B8
@82	0100F040
@83	F0001001
@84	80821000
@85	F0401882
@86	C00FF020
@87	F1A01882
@88	1882FFF8
@89	E8020008
@8A	771DF7BB
@8B	76F80000
@8C	0000003C
@8D	FFFF003A
@8E	003A76F8
@8F	F0208089
@90	0000003B
@91	76F8F6BB
@92	F7BB81D1
@93	F2740020
@94	F073F6BB
@95	4A074A06
@96	68F84000
@97	6BF88201
@98	400070E2
@99	8A128A06
@9A	000768F8
@9B	F495FFFC
@9C	018310F8
@9D	4811823A
@9E	F4E3FFFF
@9F	10F88241
@A0	018110F8
@A1	824DF073
@A2	08F8E820
@A3	826FF273
@A4	80F80001
@A5	E800F4E3
@A6	6BF80080
@A7	F6B9F7BE
@A8	0001F100
@A9	829AF073
@AA	00F87E92
@AB	6C890001
@AC	F84D0001
@AD	4E0282B2
@AE	6B0382B0
@AF	FC008222
@B0	01600001
@B1	00010000
@B2	4A074A06
@B3	00127104
@B4	8020FA4D
@B5	E5986DBB
@B6	6DEA6DBB
@B7	8030FA42
@B8	6DEA6DBB
@B9	8A07EE01
@BA	F495F6EB
@BB	F495F6EB
@BC	F495F6EB
@BD	F495F6EB
@BE	F495F6EB
@BF	F495F6EB
@C0	F495F6EB
@C1	F495F6EB
@C2	F495F6EB
@C3	81E8F273
@C4	F495F6EB
@C5	F495F6EB
@C6	81E8F273
@C7	F495F6EB
@C8	8213F273
@C9	F495F4EB
@CA	000000C4
@CB	00000724
@CC	0010803C
@CD	007EFF80
@CE	00000000
@CF	00000000
@D0	00000000
@D1	00000000
@D2	00000000
@D3	00000000
@D4	00000000
@D5	00000000
@D6	30000060
@D7	00000000
@D8	00000000
