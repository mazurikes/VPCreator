@0	200007E8
@1	08000577
@2	00000000
@3	0800057F
@4	08000585
@5	08000585
@6	08000585
@7	08000585
@8	08000585
@9	08000585
@A	080004D5
@B	08000585
@C	F802F000
@D	F1AA4483
@E	E8BA0E09
@F	47180301
@10	C178C878
@11	600C6804
@12	BF283A10
@13	4770600B
@14	F7FF4611
@15	FFF2F7FF
@16	60884955
@17	2002D1F9
@18	6800484D
@19	0008F040
@1A	F02069C0
@1B	60C87082
@1C	483DD1F9
@1D	F000F907
@1E	493870FF
@1F	61C84931
@20	49344833
@21	60482000
@22	F64F6008
@23	618830FF
@24	60C870FF
@25	49254824
@26	F04F6048
@27	491D70FF
@28	47706188
@29	F24062C8
@2A	F2426008
@2B	60C82001
@2C	40018000
@2D	C1555555
@2E	400B8000
@2F	400E8000
@30	F4106B80
@31	BD70B903
@32	F834E006
@33	D3F64295
@34	B902BD70
@35	0B02F834
@36	BF00D3F6
@37	1C402B02
@38	2200E003
@39	48154770
@3A	48114770
@3B	480D4770
@3C	6B804608
@3D	6B804805
@3E	4901200F
@3F	30000200
@40	FEFEF7FF
@41	FFB4F7FF
@42	F8334B49
@43	FF82F7FF
@44	03C4EB03
@45	03C4EB03
@46	FFB6F7FF
@47	23E0F04F
@48	60084933
@49	482FE004
@4A	6548492F
@4B	49281C40
@4C	68004825
@4D	47706008
@4E	492002C0
@4F	B5104770
@50	D1F92B80
@51	BF006023
@52	4B04F810
@53	0380F003
@54	00004770
@55	200000B0
@56	40070000
@57	E7FE4700
@58	E7FEE7FE
@59	00004770
@5A	200003E8
@5B	F828F000
@5C	B0184685
@5D	F04F0600
@5E	46AC0107
@5F	09C0E8AC
@60	FDA5F7FF
@61	E7FEBEAB
@62	007E76F8
@63	76F8FFFF
@64	FFFF0077
@65	007276F8
@66	76F8FFFF
@67	00000067
@68	006476F8
@69	FC000000
@6A	00127100
@6B	00000006
@6C	76E20012
@6D	71000003
@6E	000476E2
@6F	00127100
@70	00000006
@71	76E20012
@72	71000007
@73	000476E2
@74	00127100
@75	FF000006
@76	76E20012
@77	7100000B
@78	000476E2
@79	00127100
@7A	FFFF0006
@7B	76E20012
@7C	71000001
@7D	000476E2
@7E	FC00EE01
@7F	F000F603
@80	00127101
@81	71010001
@82	0002F000
@83	71018082
@84	88120002
@85	F0001001
@86	80824000
@87	F3101104
@88	10018182
@89	0001F040
@8A	80F8F482
@8B	F495FF88
@8C	FFFF0001
@8D	003D76F8
@8E	003976F8
@8F	F2740000
@90	F2740028
@91	000069F8
@92	003F0185
@93	018576F8
@94	F0208000
@95	F49581D1
@96	68F84A1D
@97	FFFC001D
@98	FFFF0185
@99	70E20185
@9A	8A098A0A
@9B	69F87D3F
@9C	8A078A1D
@9D	7211F4E3
@9E	0161F000
@9F	FFFF6CE9
@A0	F4E30182
@A1	10F8F4E3
@A2	88114A11
@A3	F8460160
@A4	E801F495
@A5	70E20160
@A6	FC008A11
@A7	007F0018
@A8	F6B7F4A0
@A9	82A0F84D
@AA	00127EF8
@AB	F0000011
@AC	F7B8828F
@AD	F6B882B8
@AE	F5E3F495
@AF	F6B80001
@B0	018380F8
@B1	00010000
@B2	82BE0183
@B3	F7B8EEFF
@B4	88101005
@B5	F495881A
@B6	6DBBE558
@B7	F2720002
@B8	118A1092
@B9	48130002
@BA	FC008A06
@BB	F495F495
@BC	F495F495
@BD	F495F495
@BE	F495F495
@BF	F495F495
@C0	F495F495
@C1	F495F495
@C2	F495F495
@C3	F495F495
@C4	F495F495
@C5	F495F495
@C6	F495F495
@C7	F495F495
@C8	F495F495
@C9	F495F495
@CA	00000001
@CB	080000FC
@CC	08000118
@CD	08000B0C
@CE	08000BA4
@CF	00000000
@D0	00000000
@D1	00000000
@D2	00000000
@D3	00000000
@D4	00000000
@D5	00000000
@D6	00000000
@D7	00000000
@D8	00000000
